module tmp;
    import my_pkg::*;
    int b = 5;
    initial begin
        int c = b;
    end
endmodule