`timescale 1ns/100ps

module testbench;

    logic a, b, c, r;

    truth_table DUT(
        .a ( a ),
        .b ( b ),
        .c ( c ),
        .r ( r )
    );

    `include "generator.svh"

    // TODO:
    // Референсная таблица истинности модуля 'truth_table':
    //
    // a b c   r
    // 0 0 0 | 0
    // 0 0 1 | 1
    // 0 1 0 | 1
    // 0 1 1 | 0
    // 1 0 0 | 1
    // 1 0 1 | 1
    // 1 1 0 | 0
    // 1 1 1 | 0
    //
    // Реализуйте проверку и выясните, при каких значениях
    // значения в референсной таблице не совпадают с реальными.
    //
    // Проверку можно осуществлять каждый раз, когда запускается
    // event с именем 'ev'. Отслеживайте этот момент при помощи @.
    //
    // Прототип проверки:
    //
    // initial begin
    //     logic _r;
    //     while(1) begin
    //         <ожидание event ev>;
    //         <вычисления>
    //         if( <некоторое условие> ) begin
    //             <вывод данных>;
    //         end
    //     end
    // end
    //
    // Вывод одного из значений можно реализовать, например, так:
    //
    // $display("a: %1b", a); // где 'a' - некая переменная
    //
    // Для двух значений:
    //
    // $display("a: %1b, b: %1b", b); // где 'a', 'b' - некие переменные


    // Пишите внутри этого блока
    logic tb_r;
    initial begin
        {a, b, c, tb_r} = 4'b0;
        #1
        ->> ev;
        #9
        {a, b, c, tb_r} = 4'b0011;
        #1
        ->> ev;
        #9
        {a, b, c, tb_r} = 4'b0101;
        #1
        ->> ev;
        #9
        {a, b, c, tb_r} = 4'b0110;
        #1
        ->> ev;
        #9
        {a, b, c, tb_r} = 4'b1001;
        #1
        ->> ev;
        #9
        {a, b, c, tb_r} = 4'b1011;
        #1
        ->> ev;
        #9
        {a, b, c, tb_r} = 4'b1100;
        #1
        ->> ev;
        #9
        {a, b, c, tb_r} = 4'b1110;
        #1
        ->> ev;
    end
    initial begin
        while(1) begin
            @ev;
            if (r !== tb_r) $display("a = %b, b = %b, c = %b", a, b, c);
        end
    end

endmodule
