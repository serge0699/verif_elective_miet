`timescale 1ns/100ps

module testbench;

    logic a, b, c, r;

    truth_table DUT(
        .a ( a ),
        .b ( b ),
        .c ( c ),
        .r ( r )
    );

    `include "generator.svh"

    // TODO:
    // Референсная таблица истинности модуля 'truth_table':
    //
    // a b c   r
    // 0 0 0 | 0
    // 0 0 1 | 1
    // 0 1 0 | 1
    // 0 1 1 | 0
    // 1 0 0 | 1
    // 1 0 1 | 1
    // 1 1 0 | 0
    // 1 1 1 | 0
    //
    // Реализуйте проверку и выясните, при каких значениях
    // значения в референсной таблице не совпадают с реальными.
    //
    // Проверку можно осуществлять каждый раз, когда запускается
    // event с именем 'ev'. Отслеживайте этот момент при помощи @.
    //
    // Прототип проверки:
    //
    // initial begin
    //     logic _r;
    //     while(1) begin
    //         <ожидание event ev>;
    //         <вычисления>
    //         if( <некоторое условие> ) begin
    //             <вывод данных>;
    //         end
    //     end
    // end
    //
    // Вывод одного из значений можно реализовать, например, так:
    //
    // $display("a: %1b", a); // где 'a' - некая переменная
    //
    // Для двух значений:
    //
    // $display("a: %1b, b: %1b", b); // где 'a', 'b' - некие переменные


    // Пишите внутри этого блока
    //------------------------------------------------------------
    // Считаем СДНФ по референсной таблице: b~c+a~b+b~a~c
    initial begin
        logic _r;
        while(1) begin
            @ev
            _r = !b && c || a && !b || b && !a && !c;
            if( _r != r ) begin 
                $error("incorrect truth_table");
                $display("a:%b", a, " b:%b", b, " c:%b", c); 
            end
        end
    end
    //------------------------------------------------------------

endmodule
