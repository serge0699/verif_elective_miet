`timescale 1ns/1ps

module testbench;

    logic [7:0] a;
    logic [7:0] b;
    logic       c;

    comp DUT(
        .a   ( a   ),
        .b   ( b   ),
        .c   ( c   )
    );

    // TODO:
    // Сгенерируйте входные воздействия в соответствии
    // временной диаграммой:
    //
    //     a |<----10---->|<---------------30---------------->|
    //     b |<-----------+---20---------------->|<----40---->|
    //       |            |                      |            |
    // Время |---------> 10ns ----------------> 30ns ------> 40ns
    //
    // Встройте проверки в ваш код.

    // Пишите внутри этого блока
    //------------------------------------------------------------
    initial begin
    b = 20;
    if (c != 0) $error("BAD");
    a = 10;#10ns;
    if (c != 0) $error("BAD");
    a = 30;#20ns;
    if (c != 1) $error("BAD");
    b = 40;#10ns;
    if (c != 0) $error("BAD");
    end
    //------------------------------------------------------------

endmodule
