`timescale 1ns/100ps

module testbench;

    logic [31:0] A;
    logic [31:0] B;
    logic [31:0] C;

    sum DUT(
        .a ( A ),
        .b ( B ),
        .c ( C )
    );

    `include "checker.svh"

    initial begin

        // TODO:
        // Представьте, что для каждого входного операнда (A и B)
        // интервал всех возможных значений равномерно разбит на
        // 8 одинаковых по размеру подинтервалов:
    
        // |0....|.....|.....|.....|.....|.....|.....|..max|
        // |  0  |  1  |  2  |  3  |  4  |  5  |  6  |  7  |
    
        // Ваша задача - подать значения из каждого интервала для
        // каждого операнда.
        
        // В конце симуляции будет выведена статистика о том, какая
        // часть из требуемых значений была подана. Для оценки того,
        // значения из какого интервала не были поданы, воспользуйтесь
        // отчетом 01_sum/stats/covsummary.html (отчет сформируется
        // после завершения симуляции).

        // Не забудьте про выставление задержек через '#'!

        // Пишите внутри этого блока
        //------------------------------------------------------------
        A = 32'hFFFFFFFF; B = 32'hFFFFFFFF;   
        #1ns; A = 32'h1FFFFFFF; B =32'h1FFFFFFF;
        #1ns; A = 32'h9FDCE; B =32'hB93DA; //1 <536
        #1ns; A = 32'h256667CA; B =32'h2657E698;//2 <1072
        #1ns; A = 32'h5855203F; B =32'h5E61F65A;//3 <1608

        #1ns; A = 32'h63924596; B =32'h67D97A83;//4 < 2144


        #1ns; A = 32'h8E54BADC; B =32'h8B0D2DF6;//5 <2680
        #1ns; A = 32'hBA3248CC; B =32'hB38FD0A6;//6 <3216
        #1ns; A = 32'hD89EFF9F; B =32'h44AD5E8;//7 <3752
        //------------------------------------------------------------

        -> gen_done;

    end

endmodule
