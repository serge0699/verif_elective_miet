package my_pkg;
    int b = 10;
endpackage